-- ... ...
