-- ... ...
0_0
