.- ... ... 
0_o
